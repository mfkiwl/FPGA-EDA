library verilog;
use verilog.vl_types.all;
entity XSKZQ_vlg_vec_tst is
end XSKZQ_vlg_vec_tst;
