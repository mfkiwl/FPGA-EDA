library verilog;
use verilog.vl_types.all;
entity led_xs_vlg_vec_tst is
end led_xs_vlg_vec_tst;
