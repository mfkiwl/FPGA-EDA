library verilog;
use verilog.vl_types.all;
entity LED_XS_vlg_vec_tst is
end LED_XS_vlg_vec_tst;
