library verilog;
use verilog.vl_types.all;
entity YMQ47_vlg_vec_tst is
end YMQ47_vlg_vec_tst;
