library verilog;
use verilog.vl_types.all;
entity quling_vlg_vec_tst is
end quling_vlg_vec_tst;
