library verilog;
use verilog.vl_types.all;
entity xuanze_vlg_vec_tst is
end xuanze_vlg_vec_tst;
