library verilog;
use verilog.vl_types.all;
entity YMQ58_vlg_vec_tst is
end YMQ58_vlg_vec_tst;
