library verilog;
use verilog.vl_types.all;
entity CNT24_vlg_check_tst is
    port(
        co              : in     vl_logic;
        num             : in     vl_logic_vector(4 downto 0);
        sampler_rx      : in     vl_logic
    );
end CNT24_vlg_check_tst;
