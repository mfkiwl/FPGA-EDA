LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY CTRLS IS
  PORT(CLK: IN STD_LOGIC;      
  SEL: OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END ENTITY CTRLS;
ARCHITECTURE ART OF CTRLS IS
  SIGNAL CNT: STD_LOGIC_VECTOR(2 DOWNTO 0):="000";
  BEGIN
  PROCESS(CLK) IS
    BEGIN
    IF CLK'EVENT AND CLK='1' THEN
      IF CNT="111" THEN 
         CNT<="000";
       ELSE 
         CNT<=CNT+'1';
      END IF ;
   END IF;
  END PROCESS;
  SEL<=CNT;
END ARCHITECTURE ART;

