library verilog;
use verilog.vl_types.all;
entity CNT30_vlg_vec_tst is
end CNT30_vlg_vec_tst;
