library verilog;
use verilog.vl_types.all;
entity data_change_vlg_vec_tst is
end data_change_vlg_vec_tst;
