library verilog;
use verilog.vl_types.all;
entity youxiaozhi_vlg_vec_tst is
end youxiaozhi_vlg_vec_tst;
