library verilog;
use verilog.vl_types.all;
entity TZKZQ_vlg_vec_tst is
end TZKZQ_vlg_vec_tst;
