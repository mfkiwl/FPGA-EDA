library verilog;
use verilog.vl_types.all;
entity qiuhe_vlg_vec_tst is
end qiuhe_vlg_vec_tst;
