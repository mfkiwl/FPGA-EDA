library verilog;
use verilog.vl_types.all;
entity AD0809_vlg_vec_tst is
end AD0809_vlg_vec_tst;
