library verilog;
use verilog.vl_types.all;
entity CNT24_vlg_vec_tst is
end CNT24_vlg_vec_tst;
