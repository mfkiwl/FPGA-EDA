library verilog;
use verilog.vl_types.all;
entity quzhiliu_vlg_vec_tst is
end quzhiliu_vlg_vec_tst;
