 --DTCNT9999.VHDL
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY DTCNT9999 IS
	PORT(CLK1:IN STD_LOGIC;
		  CLR:IN STD_LOGIC;
		  ENA:IN STD_LOGIC;
		  CLK2:IN STD_LOGIC;
		  COM:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		  SEG:OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENTITY DTCNT9999;
ARCHITECTURE ART OF DTCNT9999 IS
	COMPONENT CNT10 IS
		PORT(CLK:IN STD_LOGIC;
			  CLR:IN STD_LOGIC;
			  ENA:IN STD_LOGIC;
			  CQ:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
			  CO:OUT STD_LOGIC);
	END COMPONENT CNT10;
	COMPONENT CTRLS IS
		PORT(CLK:IN STD_LOGIC;
			  SEL:OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
	END COMPONENT CTRLS;
	COMPONENT DISPLAY IS
		PORT(SEL:IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			  DATAIN:IN STD_LOGIC_VECTOR(23 DOWNTO 0);
			  COM: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			  SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
	END COMPONENT DISPLAY;	
	SIGNAL S1,S2,S3,S4,S5,S6:STD_LOGIC;
	SIGNAL S:STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL DOUT:STD_LOGIC_VECTOR(23 DOWNTO 0);
	BEGIN
	U1:CNT10  PORT MAP(CLK1,CLR,ENA,DOUT(3 DOWNTO 0),S1);
	U2:CNT10  PORT MAP(S1,CLR,ENA,DOUT(7 DOWNTO 4),S2);
	U3:CNT10  PORT MAP(S2,CLR,ENA,DOUT(11 DOWNTO 8),S3);
	U4:CNT10  PORT MAP(S3,CLR,ENA,DOUT(15 DOWNTO 12),S4);
	U5:CNT10  PORT MAP(S4,CLR,ENA,DOUT(19 DOWNTO 16),S5);
	U6:CNT10  PORT MAP(S5,CLR,ENA,DOUT(23 DOWNTO 20),S6);
	U9:CTRLS  PORT MAP(CLK2,S(2 DOWNTO 0));
	U10:DISPLAY PORT MAP(S,DOUT,COM,SEG);
END ARCHITECTURE ART;
