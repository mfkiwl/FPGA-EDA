library verilog;
use verilog.vl_types.all;
entity qiuhe_gong_vlg_vec_tst is
end qiuhe_gong_vlg_vec_tst;
