library verilog;
use verilog.vl_types.all;
entity gonglvyinsu_vlg_vec_tst is
end gonglvyinsu_vlg_vec_tst;
