library verilog;
use verilog.vl_types.all;
entity wugong_vlg_vec_tst is
end wugong_vlg_vec_tst;
