library verilog;
use verilog.vl_types.all;
entity CNT60_vlg_vec_tst is
end CNT60_vlg_vec_tst;
