library verilog;
use verilog.vl_types.all;
entity yougong_vlg_vec_tst is
end yougong_vlg_vec_tst;
