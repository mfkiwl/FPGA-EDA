library verilog;
use verilog.vl_types.all;
entity XSKZ_vlg_vec_tst is
end XSKZ_vlg_vec_tst;
