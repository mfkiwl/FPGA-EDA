library verilog;
use verilog.vl_types.all;
entity genhao_vlg_vec_tst is
end genhao_vlg_vec_tst;
