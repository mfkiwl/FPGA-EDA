library verilog;
use verilog.vl_types.all;
entity shizaigonglv_vlg_vec_tst is
end shizaigonglv_vlg_vec_tst;
