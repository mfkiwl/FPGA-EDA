library verilog;
use verilog.vl_types.all;
entity YMQ38_vlg_vec_tst is
end YMQ38_vlg_vec_tst;
