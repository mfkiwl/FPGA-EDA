library verilog;
use verilog.vl_types.all;
entity DISPLAY_vlg_vec_tst is
end DISPLAY_vlg_vec_tst;
