library verilog;
use verilog.vl_types.all;
entity CNT100_vlg_vec_tst is
end CNT100_vlg_vec_tst;
