library verilog;
use verilog.vl_types.all;
entity cnt30_vlg_vec_tst is
end cnt30_vlg_vec_tst;
