library verilog;
use verilog.vl_types.all;
entity CNT7_vlg_vec_tst is
end CNT7_vlg_vec_tst;
