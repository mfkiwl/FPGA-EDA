library verilog;
use verilog.vl_types.all;
entity fenpin_vlg_vec_tst is
end fenpin_vlg_vec_tst;
