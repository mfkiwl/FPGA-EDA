LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY DISPLAY IS
  PORT(SEL: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
       DATAIN: IN STD_LOGIC_VECTOR(23 DOWNTO 0);
       COM: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
       SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END ENTITY DISPLAY;
ARCHITECTURE ART OF DISPLAY IS
  SIGNAL DATA:STD_LOGIC_VECTOR(3 DOWNTO 0);
  BEGIN
  PROCESS(SEL) IS
    BEGIN
    CASE SEL IS
      WHEN "000" => COM<="11111110";
      WHEN "001" => COM<="11111101";
      WHEN "010" => COM<="11111011";
      WHEN "011" => COM<="11110111";
      WHEN "100" => COM<="11101111";
      WHEN "101" => COM<="11011111";
      WHEN "110" => COM<="10111111";
      WHEN "111" => COM<="01111111";
      WHEN OTHERS => COM<="11111111";
    END CASE ;
  END PROCESS;
  PROCESS(SEL) IS
    BEGIN
    CASE SEL IS
      WHEN "000" =>DATA<=DATAIN(3 DOWNTO 0);
      WHEN "001" =>DATA<=DATAIN(7 DOWNTO 4);
      WHEN "010" =>DATA<=DATAIN(11 DOWNTO 8);
      WHEN "011" =>DATA<=DATAIN(15 DOWNTO 12);
		WHEN "100" =>DATA<=DATAIN(19 DOWNTO 16);
		WHEN "101" =>DATA<=DATAIN(23 DOWNTO 20);

		
      WHEN OTHERS=>DATA<="0000";
    END CASE;
       CASE DATA IS
      WHEN "0000" => SEG<="00111111";--3FH
      WHEN "0001" => SEG<="00000110";--06H
      WHEN "0010" => SEG<="01011011";--5BH
      WHEN "0011" => SEG<="01001111";--4FH
      WHEN "0100" => SEG<="01100110";--66H
      WHEN "0101" => SEG<="01101101";--6DH
      WHEN "0110" => SEG<="01111101";--7DH
      WHEN "0111" => SEG<="00000111";--07H
      WHEN "1000" => SEG<="01111111";--7FH
      WHEN "1001" => SEG<="01101111";--6FH
      WHEN OTHERS => SEG<="00000000";--00H
   END CASE ;
 END PROCESS;
END ARCHITECTURE ART;
