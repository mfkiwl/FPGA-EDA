library verilog;
use verilog.vl_types.all;
entity CNT12_vlg_vec_tst is
end CNT12_vlg_vec_tst;
