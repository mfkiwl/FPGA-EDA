library verilog;
use verilog.vl_types.all;
entity cnt60_vlg_vec_tst is
end cnt60_vlg_vec_tst;
